// this is the first Verilog project
// goal: turn on LEDs when switches are pushed
// 07/26/2022

module proj_1 (    
    input  i_Switch_1,
    input  i_Switch_2,
    input  i_Switch_3, 
    input  i_Switch_4, 
    output o_LED_1   ,
    output o_LED_2   ,
    output o_LED_3   ,
    output o_LED_4 );

    assign o_LED_1 = i_Switch_1;
    assign o_LED_2 = i_Switch_2;
    assign o_LED_3 = i_Switch_3;
    assign o_LED_4 = i_Switch_4;


endmodule
